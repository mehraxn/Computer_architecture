
ENTITY OR2LOCAL IS
	PORT(I1, I2: IN BIT;
			O:	OUT BIT);			
END OR2LOCAL;
ARCHITECTURE gate OF OR2LOCAL IS
BEGIN	
	O <= I1 or I2;		
END gate;