
ENTITY AND2LOCAL IS
	PORT(I1, I2: IN BIT;
			O:	OUT BIT);			
END AND2LOCAL;
ARCHITECTURE gate OF AND2LOCAL IS
BEGIN	
	O <= I1 and I2;		
END gate;