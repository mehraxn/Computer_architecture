
ENTITY OR3LOCAL IS
	PORT(I1, I2, I3: IN BIT;
			O:	OUT BIT);			
END OR3LOCAL;
ARCHITECTURE gate OF OR3LOCAL IS
BEGIN	
	O <= I1 or I2 or I3;		
END gate;