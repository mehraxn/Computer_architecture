
ENTITY OR4LOCAL IS
	PORT(I1, I2, I3, I4: IN BIT;
			O:	OUT BIT);			
END OR4LOCAL;
ARCHITECTURE gate OF OR4LOCAL IS
BEGIN	
	O <= I1 or I2 or I3 or I4;		
END gate;