

ENTITY AND3LOCAL IS
	PORT(I1, I2, I3: IN BIT;
			O:	OUT BIT);			
END AND3LOCAL;
ARCHITECTURE gate OF AND3LOCAL IS
BEGIN	
	O <= I1 and I2 and I3;		
END gate;